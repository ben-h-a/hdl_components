module tb;

    

    sp_ram #(
        .WIDTH(8),
        .DEPTH(8),
        .STRB_WIDTH(8)
    ) 
    u_ram(

    );

endmodule